library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Decoder5to32 is
Port( input : in std_logic_vector( 4 downto 0);
		output : out std_logic_vector ( 31 downto 0)
		);
end Decoder5to32;

architecture Behavioral of Decoder5to32 is
signal temp_output:std_logic_vector ( 31 downto 0);

begin
temp_output<= "00000000000000000000000000000000" when input = "00000" else
		"00000000000000000000000000000010" when input = "00001" else
		"00000000000000000000000000000100" when input = "00010" else
		"00000000000000000000000000001000" when input = "00011" else
		"00000000000000000000000000010000" when input = "00100" else
		"00000000000000000000000000100000" when input = "00101" else
		"00000000000000000000000001000000" when input = "00110" else
		"00000000000000000000000010000000" when input = "00111" else
		"00000000000000000000000100000000" when input = "01000" else
		"00000000000000000000001000000000" when input = "01001" else
		"00000000000000000000010000000000" when input = "01010" else
		"00000000000000000000100000000000" when input = "01011" else
		"00000000000000000001000000000000" when input = "01100" else
		"00000000000000000010000000000000" when input = "01101" else
		"00000000000000000100000000000000" when input = "01110" else
		"00000000000000001000000000000000" when input = "01111" else
		"00000000000000010000000000000000" when input = "10000" else
		"00000000000000100000000000000000" when input = "10001" else
		"00000000000001000000000000000000" when input = "10010" else
		"00000000000010000000000000000000" when input = "10011" else
		"00000000000100000000000000000000" when input = "10100" else
		"00000000001000000000000000000000" when input = "10101" else
		"00000000010000000000000000000000" when input = "10110" else
		"00000000100000000000000000000000" when input = "10111" else
		"00000001000000000000000000000000" when input = "11000" else
		"00000010000000000000000000000000" when input = "11001" else
		"00000100000000000000000000000000" when input = "11010" else
		"00001000000000000000000000000000" when input = "11011" else
		"00010000000000000000000000000000" when input = "11100" else
		"00100000000000000000000000000000" when input = "11101" else
		"01000000000000000000000000000000" when input = "11110" else
		"10000000000000000000000000000000" when input = "11111";
		
		output<=temp_output after 5 ns;



end Behavioral;