library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity CONTROL is
end CONTROL;

architecture Behavioral of CONTROL is

begin


end Behavioral;

